`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.02.2019 18:36:19
// Design Name: 
// Module Name: Sig_ROM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Sig_ROM(
    input           clk,
    input   [9:0]   x,
    output  [15:0]  out
    );
    
    reg [15:0] mem [1023:0];
    reg [9:0] y;
    
    always @(posedge clk)
    begin
        if($signed(x) >= 0)
            y <= x+512;
        else 
            y <= x-512;      
    end
        
    initial
    begin
    mem[ 0 ] = 16'b0000000000001010;
    mem[ 1 ] = 16'b0000000000001011;
    mem[ 2 ] = 16'b0000000000001011;
    mem[ 3 ] = 16'b0000000000001011;
    mem[ 4 ] = 16'b0000000000001011;
    mem[ 5 ] = 16'b0000000000001011;
    mem[ 6 ] = 16'b0000000000001100;
    mem[ 7 ] = 16'b0000000000001100;
    mem[ 8 ] = 16'b0000000000001100;
    mem[ 9 ] = 16'b0000000000001100;
    mem[ 10 ] = 16'b0000000000001100;
    mem[ 11 ] = 16'b0000000000001101;
    mem[ 12 ] = 16'b0000000000001101;
    mem[ 13 ] = 16'b0000000000001101;
    mem[ 14 ] = 16'b0000000000001101;
    mem[ 15 ] = 16'b0000000000001101;
    mem[ 16 ] = 16'b0000000000001110;
    mem[ 17 ] = 16'b0000000000001110;
    mem[ 18 ] = 16'b0000000000001110;
    mem[ 19 ] = 16'b0000000000001110;
    mem[ 20 ] = 16'b0000000000001111;
    mem[ 21 ] = 16'b0000000000001111;
    mem[ 22 ] = 16'b0000000000001111;
    mem[ 23 ] = 16'b0000000000001111;
    mem[ 24 ] = 16'b0000000000001111;
    mem[ 25 ] = 16'b0000000000010000;
    mem[ 26 ] = 16'b0000000000010000;
    mem[ 27 ] = 16'b0000000000010000;
    mem[ 28 ] = 16'b0000000000010001;
    mem[ 29 ] = 16'b0000000000010001;
    mem[ 30 ] = 16'b0000000000010001;
    mem[ 31 ] = 16'b0000000000010001;
    mem[ 32 ] = 16'b0000000000010010;
    mem[ 33 ] = 16'b0000000000010010;
    mem[ 34 ] = 16'b0000000000010010;
    mem[ 35 ] = 16'b0000000000010010;
    mem[ 36 ] = 16'b0000000000010011;
    mem[ 37 ] = 16'b0000000000010011;
    mem[ 38 ] = 16'b0000000000010011;
    mem[ 39 ] = 16'b0000000000010100;
    mem[ 40 ] = 16'b0000000000010100;
    mem[ 41 ] = 16'b0000000000010100;
    mem[ 42 ] = 16'b0000000000010101;
    mem[ 43 ] = 16'b0000000000010101;
    mem[ 44 ] = 16'b0000000000010101;
    mem[ 45 ] = 16'b0000000000010110;
    mem[ 46 ] = 16'b0000000000010110;
    mem[ 47 ] = 16'b0000000000010110;
    mem[ 48 ] = 16'b0000000000010111;
    mem[ 49 ] = 16'b0000000000010111;
    mem[ 50 ] = 16'b0000000000010111;
    mem[ 51 ] = 16'b0000000000011000;
    mem[ 52 ] = 16'b0000000000011000;
    mem[ 53 ] = 16'b0000000000011001;
    mem[ 54 ] = 16'b0000000000011001;
    mem[ 55 ] = 16'b0000000000011001;
    mem[ 56 ] = 16'b0000000000011010;
    mem[ 57 ] = 16'b0000000000011010;
    mem[ 58 ] = 16'b0000000000011011;
    mem[ 59 ] = 16'b0000000000011011;
    mem[ 60 ] = 16'b0000000000011100;
    mem[ 61 ] = 16'b0000000000011100;
    mem[ 62 ] = 16'b0000000000011100;
    mem[ 63 ] = 16'b0000000000011101;
    mem[ 64 ] = 16'b0000000000011101;
    mem[ 65 ] = 16'b0000000000011110;
    mem[ 66 ] = 16'b0000000000011110;
    mem[ 67 ] = 16'b0000000000011111;
    mem[ 68 ] = 16'b0000000000011111;
    mem[ 69 ] = 16'b0000000000100000;
    mem[ 70 ] = 16'b0000000000100000;
    mem[ 71 ] = 16'b0000000000100001;
    mem[ 72 ] = 16'b0000000000100001;
    mem[ 73 ] = 16'b0000000000100010;
    mem[ 74 ] = 16'b0000000000100010;
    mem[ 75 ] = 16'b0000000000100011;
    mem[ 76 ] = 16'b0000000000100100;
    mem[ 77 ] = 16'b0000000000100100;
    mem[ 78 ] = 16'b0000000000100101;
    mem[ 79 ] = 16'b0000000000100101;
    mem[ 80 ] = 16'b0000000000100110;
    mem[ 81 ] = 16'b0000000000100110;
    mem[ 82 ] = 16'b0000000000100111;
    mem[ 83 ] = 16'b0000000000101000;
    mem[ 84 ] = 16'b0000000000101000;
    mem[ 85 ] = 16'b0000000000101001;
    mem[ 86 ] = 16'b0000000000101010;
    mem[ 87 ] = 16'b0000000000101010;
    mem[ 88 ] = 16'b0000000000101011;
    mem[ 89 ] = 16'b0000000000101100;
    mem[ 90 ] = 16'b0000000000101100;
    mem[ 91 ] = 16'b0000000000101101;
    mem[ 92 ] = 16'b0000000000101110;
    mem[ 93 ] = 16'b0000000000101110;
    mem[ 94 ] = 16'b0000000000101111;
    mem[ 95 ] = 16'b0000000000110000;
    mem[ 96 ] = 16'b0000000000110001;
    mem[ 97 ] = 16'b0000000000110001;
    mem[ 98 ] = 16'b0000000000110010;
    mem[ 99 ] = 16'b0000000000110011;
    mem[ 100 ] = 16'b0000000000110100;
    mem[ 101 ] = 16'b0000000000110101;
    mem[ 102 ] = 16'b0000000000110110;
    mem[ 103 ] = 16'b0000000000110110;
    mem[ 104 ] = 16'b0000000000110111;
    mem[ 105 ] = 16'b0000000000111000;
    mem[ 106 ] = 16'b0000000000111001;
    mem[ 107 ] = 16'b0000000000111010;
    mem[ 108 ] = 16'b0000000000111011;
    mem[ 109 ] = 16'b0000000000111100;
    mem[ 110 ] = 16'b0000000000111101;
    mem[ 111 ] = 16'b0000000000111110;
    mem[ 112 ] = 16'b0000000000111111;
    mem[ 113 ] = 16'b0000000001000000;
    mem[ 114 ] = 16'b0000000001000001;
    mem[ 115 ] = 16'b0000000001000010;
    mem[ 116 ] = 16'b0000000001000011;
    mem[ 117 ] = 16'b0000000001000100;
    mem[ 118 ] = 16'b0000000001000101;
    mem[ 119 ] = 16'b0000000001000110;
    mem[ 120 ] = 16'b0000000001000111;
    mem[ 121 ] = 16'b0000000001001000;
    mem[ 122 ] = 16'b0000000001001001;
    mem[ 123 ] = 16'b0000000001001010;
    mem[ 124 ] = 16'b0000000001001100;
    mem[ 125 ] = 16'b0000000001001101;
    mem[ 126 ] = 16'b0000000001001110;
    mem[ 127 ] = 16'b0000000001001111;
    mem[ 128 ] = 16'b0000000001010001;
    mem[ 129 ] = 16'b0000000001010010;
    mem[ 130 ] = 16'b0000000001010011;
    mem[ 131 ] = 16'b0000000001010100;
    mem[ 132 ] = 16'b0000000001010110;
    mem[ 133 ] = 16'b0000000001010111;
    mem[ 134 ] = 16'b0000000001011000;
    mem[ 135 ] = 16'b0000000001011010;
    mem[ 136 ] = 16'b0000000001011011;
    mem[ 137 ] = 16'b0000000001011101;
    mem[ 138 ] = 16'b0000000001011110;
    mem[ 139 ] = 16'b0000000001100000;
    mem[ 140 ] = 16'b0000000001100001;
    mem[ 141 ] = 16'b0000000001100011;
    mem[ 142 ] = 16'b0000000001100100;
    mem[ 143 ] = 16'b0000000001100110;
    mem[ 144 ] = 16'b0000000001100111;
    mem[ 145 ] = 16'b0000000001101001;
    mem[ 146 ] = 16'b0000000001101011;
    mem[ 147 ] = 16'b0000000001101100;
    mem[ 148 ] = 16'b0000000001101110;
    mem[ 149 ] = 16'b0000000001110000;
    mem[ 150 ] = 16'b0000000001110010;
    mem[ 151 ] = 16'b0000000001110011;
    mem[ 152 ] = 16'b0000000001110101;
    mem[ 153 ] = 16'b0000000001110111;
    mem[ 154 ] = 16'b0000000001111001;
    mem[ 155 ] = 16'b0000000001111011;
    mem[ 156 ] = 16'b0000000001111101;
    mem[ 157 ] = 16'b0000000001111111;
    mem[ 158 ] = 16'b0000000010000001;
    mem[ 159 ] = 16'b0000000010000011;
    mem[ 160 ] = 16'b0000000010000101;
    mem[ 161 ] = 16'b0000000010000111;
    mem[ 162 ] = 16'b0000000010001001;
    mem[ 163 ] = 16'b0000000010001011;
    mem[ 164 ] = 16'b0000000010001101;
    mem[ 165 ] = 16'b0000000010010000;
    mem[ 166 ] = 16'b0000000010010010;
    mem[ 167 ] = 16'b0000000010010100;
    mem[ 168 ] = 16'b0000000010010111;
    mem[ 169 ] = 16'b0000000010011001;
    mem[ 170 ] = 16'b0000000010011011;
    mem[ 171 ] = 16'b0000000010011110;
    mem[ 172 ] = 16'b0000000010100000;
    mem[ 173 ] = 16'b0000000010100011;
    mem[ 174 ] = 16'b0000000010100101;
    mem[ 175 ] = 16'b0000000010101000;
    mem[ 176 ] = 16'b0000000010101011;
    mem[ 177 ] = 16'b0000000010101101;
    mem[ 178 ] = 16'b0000000010110000;
    mem[ 179 ] = 16'b0000000010110011;
    mem[ 180 ] = 16'b0000000010110110;
    mem[ 181 ] = 16'b0000000010111000;
    mem[ 182 ] = 16'b0000000010111011;
    mem[ 183 ] = 16'b0000000010111110;
    mem[ 184 ] = 16'b0000000011000001;
    mem[ 185 ] = 16'b0000000011000100;
    mem[ 186 ] = 16'b0000000011000111;
    mem[ 187 ] = 16'b0000000011001010;
    mem[ 188 ] = 16'b0000000011001110;
    mem[ 189 ] = 16'b0000000011010001;
    mem[ 190 ] = 16'b0000000011010100;
    mem[ 191 ] = 16'b0000000011010111;
    mem[ 192 ] = 16'b0000000011011011;
    mem[ 193 ] = 16'b0000000011011110;
    mem[ 194 ] = 16'b0000000011100010;
    mem[ 195 ] = 16'b0000000011100101;
    mem[ 196 ] = 16'b0000000011101001;
    mem[ 197 ] = 16'b0000000011101101;
    mem[ 198 ] = 16'b0000000011110000;
    mem[ 199 ] = 16'b0000000011110100;
    mem[ 200 ] = 16'b0000000011111000;
    mem[ 201 ] = 16'b0000000011111100;
    mem[ 202 ] = 16'b0000000100000000;
    mem[ 203 ] = 16'b0000000100000100;
    mem[ 204 ] = 16'b0000000100001000;
    mem[ 205 ] = 16'b0000000100001100;
    mem[ 206 ] = 16'b0000000100010000;
    mem[ 207 ] = 16'b0000000100010100;
    mem[ 208 ] = 16'b0000000100011001;
    mem[ 209 ] = 16'b0000000100011101;
    mem[ 210 ] = 16'b0000000100100001;
    mem[ 211 ] = 16'b0000000100100110;
    mem[ 212 ] = 16'b0000000100101011;
    mem[ 213 ] = 16'b0000000100101111;
    mem[ 214 ] = 16'b0000000100110100;
    mem[ 215 ] = 16'b0000000100111001;
    mem[ 216 ] = 16'b0000000100111110;
    mem[ 217 ] = 16'b0000000101000011;
    mem[ 218 ] = 16'b0000000101001000;
    mem[ 219 ] = 16'b0000000101001101;
    mem[ 220 ] = 16'b0000000101010010;
    mem[ 221 ] = 16'b0000000101010111;
    mem[ 222 ] = 16'b0000000101011101;
    mem[ 223 ] = 16'b0000000101100010;
    mem[ 224 ] = 16'b0000000101101000;
    mem[ 225 ] = 16'b0000000101101101;
    mem[ 226 ] = 16'b0000000101110011;
    mem[ 227 ] = 16'b0000000101111001;
    mem[ 228 ] = 16'b0000000101111110;
    mem[ 229 ] = 16'b0000000110000100;
    mem[ 230 ] = 16'b0000000110001010;
    mem[ 231 ] = 16'b0000000110010001;
    mem[ 232 ] = 16'b0000000110010111;
    mem[ 233 ] = 16'b0000000110011101;
    mem[ 234 ] = 16'b0000000110100100;
    mem[ 235 ] = 16'b0000000110101010;
    mem[ 236 ] = 16'b0000000110110001;
    mem[ 237 ] = 16'b0000000110111000;
    mem[ 238 ] = 16'b0000000110111110;
    mem[ 239 ] = 16'b0000000111000101;
    mem[ 240 ] = 16'b0000000111001100;
    mem[ 241 ] = 16'b0000000111010011;
    mem[ 242 ] = 16'b0000000111011011;
    mem[ 243 ] = 16'b0000000111100010;
    mem[ 244 ] = 16'b0000000111101010;
    mem[ 245 ] = 16'b0000000111110001;
    mem[ 246 ] = 16'b0000000111111001;
    mem[ 247 ] = 16'b0000001000000001;
    mem[ 248 ] = 16'b0000001000001001;
    mem[ 249 ] = 16'b0000001000010001;
    mem[ 250 ] = 16'b0000001000011001;
    mem[ 251 ] = 16'b0000001000100001;
    mem[ 252 ] = 16'b0000001000101010;
    mem[ 253 ] = 16'b0000001000110010;
    mem[ 254 ] = 16'b0000001000111011;
    mem[ 255 ] = 16'b0000001001000100;
    mem[ 256 ] = 16'b0000001001001101;
    mem[ 257 ] = 16'b0000001001010110;
    mem[ 258 ] = 16'b0000001001011111;
    mem[ 259 ] = 16'b0000001001101001;
    mem[ 260 ] = 16'b0000001001110010;
    mem[ 261 ] = 16'b0000001001111100;
    mem[ 262 ] = 16'b0000001010000110;
    mem[ 263 ] = 16'b0000001010010000;
    mem[ 264 ] = 16'b0000001010011010;
    mem[ 265 ] = 16'b0000001010100100;
    mem[ 266 ] = 16'b0000001010101110;
    mem[ 267 ] = 16'b0000001010111001;
    mem[ 268 ] = 16'b0000001011000100;
    mem[ 269 ] = 16'b0000001011001111;
    mem[ 270 ] = 16'b0000001011011010;
    mem[ 271 ] = 16'b0000001011100101;
    mem[ 272 ] = 16'b0000001011110000;
    mem[ 273 ] = 16'b0000001011111100;
    mem[ 274 ] = 16'b0000001100001000;
    mem[ 275 ] = 16'b0000001100010100;
    mem[ 276 ] = 16'b0000001100100000;
    mem[ 277 ] = 16'b0000001100101100;
    mem[ 278 ] = 16'b0000001100111001;
    mem[ 279 ] = 16'b0000001101000101;
    mem[ 280 ] = 16'b0000001101010010;
    mem[ 281 ] = 16'b0000001101011111;
    mem[ 282 ] = 16'b0000001101101100;
    mem[ 283 ] = 16'b0000001101111010;
    mem[ 284 ] = 16'b0000001110000111;
    mem[ 285 ] = 16'b0000001110010101;
    mem[ 286 ] = 16'b0000001110100011;
    mem[ 287 ] = 16'b0000001110110010;
    mem[ 288 ] = 16'b0000001111000000;
    mem[ 289 ] = 16'b0000001111001111;
    mem[ 290 ] = 16'b0000001111011110;
    mem[ 291 ] = 16'b0000001111101101;
    mem[ 292 ] = 16'b0000001111111100;
    mem[ 293 ] = 16'b0000010000001100;
    mem[ 294 ] = 16'b0000010000011011;
    mem[ 295 ] = 16'b0000010000101011;
    mem[ 296 ] = 16'b0000010000111100;
    mem[ 297 ] = 16'b0000010001001100;
    mem[ 298 ] = 16'b0000010001011101;
    mem[ 299 ] = 16'b0000010001101110;
    mem[ 300 ] = 16'b0000010001111111;
    mem[ 301 ] = 16'b0000010010010001;
    mem[ 302 ] = 16'b0000010010100010;
    mem[ 303 ] = 16'b0000010010110100;
    mem[ 304 ] = 16'b0000010011000111;
    mem[ 305 ] = 16'b0000010011011001;
    mem[ 306 ] = 16'b0000010011101100;
    mem[ 307 ] = 16'b0000010011111111;
    mem[ 308 ] = 16'b0000010100010010;
    mem[ 309 ] = 16'b0000010100100110;
    mem[ 310 ] = 16'b0000010100111010;
    mem[ 311 ] = 16'b0000010101001110;
    mem[ 312 ] = 16'b0000010101100011;
    mem[ 313 ] = 16'b0000010101110111;
    mem[ 314 ] = 16'b0000010110001101;
    mem[ 315 ] = 16'b0000010110100010;
    mem[ 316 ] = 16'b0000010110111000;
    mem[ 317 ] = 16'b0000010111001110;
    mem[ 318 ] = 16'b0000010111100100;
    mem[ 319 ] = 16'b0000010111111011;
    mem[ 320 ] = 16'b0000011000010010;
    mem[ 321 ] = 16'b0000011000101001;
    mem[ 322 ] = 16'b0000011001000000;
    mem[ 323 ] = 16'b0000011001011000;
    mem[ 324 ] = 16'b0000011001110001;
    mem[ 325 ] = 16'b0000011010001001;
    mem[ 326 ] = 16'b0000011010100010;
    mem[ 327 ] = 16'b0000011010111100;
    mem[ 328 ] = 16'b0000011011010101;
    mem[ 329 ] = 16'b0000011011101111;
    mem[ 330 ] = 16'b0000011100001010;
    mem[ 331 ] = 16'b0000011100100101;
    mem[ 332 ] = 16'b0000011101000000;
    mem[ 333 ] = 16'b0000011101011011;
    mem[ 334 ] = 16'b0000011101110111;
    mem[ 335 ] = 16'b0000011110010100;
    mem[ 336 ] = 16'b0000011110110000;
    mem[ 337 ] = 16'b0000011111001110;
    mem[ 338 ] = 16'b0000011111101011;
    mem[ 339 ] = 16'b0000100000001001;
    mem[ 340 ] = 16'b0000100000100111;
    mem[ 341 ] = 16'b0000100001000110;
    mem[ 342 ] = 16'b0000100001100101;
    mem[ 343 ] = 16'b0000100010000101;
    mem[ 344 ] = 16'b0000100010100101;
    mem[ 345 ] = 16'b0000100011000101;
    mem[ 346 ] = 16'b0000100011100110;
    mem[ 347 ] = 16'b0000100100001000;
    mem[ 348 ] = 16'b0000100100101001;
    mem[ 349 ] = 16'b0000100101001100;
    mem[ 350 ] = 16'b0000100101101110;
    mem[ 351 ] = 16'b0000100110010010;
    mem[ 352 ] = 16'b0000100110110101;
    mem[ 353 ] = 16'b0000100111011001;
    mem[ 354 ] = 16'b0000100111111110;
    mem[ 355 ] = 16'b0000101000100011;
    mem[ 356 ] = 16'b0000101001001001;
    mem[ 357 ] = 16'b0000101001101111;
    mem[ 358 ] = 16'b0000101010010101;
    mem[ 359 ] = 16'b0000101010111100;
    mem[ 360 ] = 16'b0000101011100100;
    mem[ 361 ] = 16'b0000101100001100;
    mem[ 362 ] = 16'b0000101100110101;
    mem[ 363 ] = 16'b0000101101011110;
    mem[ 364 ] = 16'b0000101110001000;
    mem[ 365 ] = 16'b0000101110110010;
    mem[ 366 ] = 16'b0000101111011101;
    mem[ 367 ] = 16'b0000110000001000;
    mem[ 368 ] = 16'b0000110000110100;
    mem[ 369 ] = 16'b0000110001100000;
    mem[ 370 ] = 16'b0000110010001101;
    mem[ 371 ] = 16'b0000110010111011;
    mem[ 372 ] = 16'b0000110011101001;
    mem[ 373 ] = 16'b0000110100011000;
    mem[ 374 ] = 16'b0000110101000111;
    mem[ 375 ] = 16'b0000110101110111;
    mem[ 376 ] = 16'b0000110110101000;
    mem[ 377 ] = 16'b0000110111011001;
    mem[ 378 ] = 16'b0000111000001010;
    mem[ 379 ] = 16'b0000111000111101;
    mem[ 380 ] = 16'b0000111001110000;
    mem[ 381 ] = 16'b0000111010100011;
    mem[ 382 ] = 16'b0000111011010111;
    mem[ 383 ] = 16'b0000111100001100;
    mem[ 384 ] = 16'b0000111101000010;
    mem[ 385 ] = 16'b0000111101111000;
    mem[ 386 ] = 16'b0000111110101110;
    mem[ 387 ] = 16'b0000111111100110;
    mem[ 388 ] = 16'b0001000000011110;
    mem[ 389 ] = 16'b0001000001010110;
    mem[ 390 ] = 16'b0001000010010000;
    mem[ 391 ] = 16'b0001000011001010;
    mem[ 392 ] = 16'b0001000100000100;
    mem[ 393 ] = 16'b0001000101000000;
    mem[ 394 ] = 16'b0001000101111100;
    mem[ 395 ] = 16'b0001000110111001;
    mem[ 396 ] = 16'b0001000111110110;
    mem[ 397 ] = 16'b0001001000110100;
    mem[ 398 ] = 16'b0001001001110011;
    mem[ 399 ] = 16'b0001001010110010;
    mem[ 400 ] = 16'b0001001011110011;
    mem[ 401 ] = 16'b0001001100110100;
    mem[ 402 ] = 16'b0001001101110101;
    mem[ 403 ] = 16'b0001001110111000;
    mem[ 404 ] = 16'b0001001111111011;
    mem[ 405 ] = 16'b0001010000111111;
    mem[ 406 ] = 16'b0001010010000011;
    mem[ 407 ] = 16'b0001010011001000;
    mem[ 408 ] = 16'b0001010100001110;
    mem[ 409 ] = 16'b0001010101010101;
    mem[ 410 ] = 16'b0001010110011101;
    mem[ 411 ] = 16'b0001010111100101;
    mem[ 412 ] = 16'b0001011000101110;
    mem[ 413 ] = 16'b0001011001111000;
    mem[ 414 ] = 16'b0001011011000010;
    mem[ 415 ] = 16'b0001011100001101;
    mem[ 416 ] = 16'b0001011101011001;
    mem[ 417 ] = 16'b0001011110100110;
    mem[ 418 ] = 16'b0001011111110011;
    mem[ 419 ] = 16'b0001100001000010;
    mem[ 420 ] = 16'b0001100010010001;
    mem[ 421 ] = 16'b0001100011100001;
    mem[ 422 ] = 16'b0001100100110001;
    mem[ 423 ] = 16'b0001100110000010;
    mem[ 424 ] = 16'b0001100111010101;
    mem[ 425 ] = 16'b0001101000100111;
    mem[ 426 ] = 16'b0001101001111011;
    mem[ 427 ] = 16'b0001101011001111;
    mem[ 428 ] = 16'b0001101100100101;
    mem[ 429 ] = 16'b0001101101111011;
    mem[ 430 ] = 16'b0001101111010001;
    mem[ 431 ] = 16'b0001110000101001;
    mem[ 432 ] = 16'b0001110010000001;
    mem[ 433 ] = 16'b0001110011011010;
    mem[ 434 ] = 16'b0001110100110100;
    mem[ 435 ] = 16'b0001110110001110;
    mem[ 436 ] = 16'b0001110111101010;
    mem[ 437 ] = 16'b0001111001000110;
    mem[ 438 ] = 16'b0001111010100010;
    mem[ 439 ] = 16'b0001111100000000;
    mem[ 440 ] = 16'b0001111101011110;
    mem[ 441 ] = 16'b0001111110111110;
    mem[ 442 ] = 16'b0010000000011101;
    mem[ 443 ] = 16'b0010000001111110;
    mem[ 444 ] = 16'b0010000011011111;
    mem[ 445 ] = 16'b0010000101000001;
    mem[ 446 ] = 16'b0010000110100100;
    mem[ 447 ] = 16'b0010001000001000;
    mem[ 448 ] = 16'b0010001001101100;
    mem[ 449 ] = 16'b0010001011010001;
    mem[ 450 ] = 16'b0010001100110111;
    mem[ 451 ] = 16'b0010001110011101;
    mem[ 452 ] = 16'b0010010000000101;
    mem[ 453 ] = 16'b0010010001101100;
    mem[ 454 ] = 16'b0010010011010101;
    mem[ 455 ] = 16'b0010010100111110;
    mem[ 456 ] = 16'b0010010110101000;
    mem[ 457 ] = 16'b0010011000010011;
    mem[ 458 ] = 16'b0010011001111110;
    mem[ 459 ] = 16'b0010011011101010;
    mem[ 460 ] = 16'b0010011101010111;
    mem[ 461 ] = 16'b0010011111000100;
    mem[ 462 ] = 16'b0010100000110010;
    mem[ 463 ] = 16'b0010100010100001;
    mem[ 464 ] = 16'b0010100100010000;
    mem[ 465 ] = 16'b0010100110000000;
    mem[ 466 ] = 16'b0010100111110001;
    mem[ 467 ] = 16'b0010101001100010;
    mem[ 468 ] = 16'b0010101011010011;
    mem[ 469 ] = 16'b0010101101000110;
    mem[ 470 ] = 16'b0010101110111000;
    mem[ 471 ] = 16'b0010110000101100;
    mem[ 472 ] = 16'b0010110010100000;
    mem[ 473 ] = 16'b0010110100010100;
    mem[ 474 ] = 16'b0010110110001010;
    mem[ 475 ] = 16'b0010110111111111;
    mem[ 476 ] = 16'b0010111001110101;
    mem[ 477 ] = 16'b0010111011101100;
    mem[ 478 ] = 16'b0010111101100011;
    mem[ 479 ] = 16'b0010111111011011;
    mem[ 480 ] = 16'b0011000001010011;
    mem[ 481 ] = 16'b0011000011001011;
    mem[ 482 ] = 16'b0011000101000100;
    mem[ 483 ] = 16'b0011000110111110;
    mem[ 484 ] = 16'b0011001000111000;
    mem[ 485 ] = 16'b0011001010110010;
    mem[ 486 ] = 16'b0011001100101101;
    mem[ 487 ] = 16'b0011001110101000;
    mem[ 488 ] = 16'b0011010000100011;
    mem[ 489 ] = 16'b0011010010011111;
    mem[ 490 ] = 16'b0011010100011011;
    mem[ 491 ] = 16'b0011010110010111;
    mem[ 492 ] = 16'b0011011000010100;
    mem[ 493 ] = 16'b0011011010010001;
    mem[ 494 ] = 16'b0011011100001111;
    mem[ 495 ] = 16'b0011011110001100;
    mem[ 496 ] = 16'b0011100000001010;
    mem[ 497 ] = 16'b0011100010001000;
    mem[ 498 ] = 16'b0011100100000111;
    mem[ 499 ] = 16'b0011100110000101;
    mem[ 500 ] = 16'b0011101000000100;
    mem[ 501 ] = 16'b0011101010000011;
    mem[ 502 ] = 16'b0011101100000010;
    mem[ 503 ] = 16'b0011101110000001;
    mem[ 504 ] = 16'b0011110000000001;
    mem[ 505 ] = 16'b0011110010000000;
    mem[ 506 ] = 16'b0011110100000000;
    mem[ 507 ] = 16'b0011110110000000;
    mem[ 508 ] = 16'b0011111000000000;
    mem[ 509 ] = 16'b0011111010000000;
    mem[ 510 ] = 16'b0011111100000000;
    mem[ 511 ] = 16'b0011111110000000;
    mem[ 512 ] = 16'b0100000000000000;
    mem[ 513 ] = 16'b0100000001111111;
    mem[ 514 ] = 16'b0100000011111111;
    mem[ 515 ] = 16'b0100000101111111;
    mem[ 516 ] = 16'b0100000111111111;
    mem[ 517 ] = 16'b0100001001111111;
    mem[ 518 ] = 16'b0100001011111111;
    mem[ 519 ] = 16'b0100001101111111;
    mem[ 520 ] = 16'b0100001111111110;
    mem[ 521 ] = 16'b0100010001111110;
    mem[ 522 ] = 16'b0100010011111101;
    mem[ 523 ] = 16'b0100010101111100;
    mem[ 524 ] = 16'b0100010111111011;
    mem[ 525 ] = 16'b0100011001111010;
    mem[ 526 ] = 16'b0100011011111000;
    mem[ 527 ] = 16'b0100011101110111;
    mem[ 528 ] = 16'b0100011111110101;
    mem[ 529 ] = 16'b0100100001110011;
    mem[ 530 ] = 16'b0100100011110000;
    mem[ 531 ] = 16'b0100100101101110;
    mem[ 532 ] = 16'b0100100111101011;
    mem[ 533 ] = 16'b0100101001101000;
    mem[ 534 ] = 16'b0100101011100100;
    mem[ 535 ] = 16'b0100101101100000;
    mem[ 536 ] = 16'b0100101111011100;
    mem[ 537 ] = 16'b0100110001010111;
    mem[ 538 ] = 16'b0100110011010010;
    mem[ 539 ] = 16'b0100110101001101;
    mem[ 540 ] = 16'b0100110111000111;
    mem[ 541 ] = 16'b0100111001000001;
    mem[ 542 ] = 16'b0100111010111011;
    mem[ 543 ] = 16'b0100111100110100;
    mem[ 544 ] = 16'b0100111110101100;
    mem[ 545 ] = 16'b0101000000100100;
    mem[ 546 ] = 16'b0101000010011100;
    mem[ 547 ] = 16'b0101000100010011;
    mem[ 548 ] = 16'b0101000110001010;
    mem[ 549 ] = 16'b0101001000000000;
    mem[ 550 ] = 16'b0101001001110101;
    mem[ 551 ] = 16'b0101001011101011;
    mem[ 552 ] = 16'b0101001101011111;
    mem[ 553 ] = 16'b0101001111010011;
    mem[ 554 ] = 16'b0101010001000111;
    mem[ 555 ] = 16'b0101010010111001;
    mem[ 556 ] = 16'b0101010100101100;
    mem[ 557 ] = 16'b0101010110011101;
    mem[ 558 ] = 16'b0101011000001110;
    mem[ 559 ] = 16'b0101011001111111;
    mem[ 560 ] = 16'b0101011011101111;
    mem[ 561 ] = 16'b0101011101011110;
    mem[ 562 ] = 16'b0101011111001101;
    mem[ 563 ] = 16'b0101100000111011;
    mem[ 564 ] = 16'b0101100010101000;
    mem[ 565 ] = 16'b0101100100010101;
    mem[ 566 ] = 16'b0101100110000001;
    mem[ 567 ] = 16'b0101100111101100;
    mem[ 568 ] = 16'b0101101001010111;
    mem[ 569 ] = 16'b0101101011000001;
    mem[ 570 ] = 16'b0101101100101010;
    mem[ 571 ] = 16'b0101101110010011;
    mem[ 572 ] = 16'b0101101111111010;
    mem[ 573 ] = 16'b0101110001100010;
    mem[ 574 ] = 16'b0101110011001000;
    mem[ 575 ] = 16'b0101110100101110;
    mem[ 576 ] = 16'b0101110110010011;
    mem[ 577 ] = 16'b0101110111110111;
    mem[ 578 ] = 16'b0101111001011011;
    mem[ 579 ] = 16'b0101111010111110;
    mem[ 580 ] = 16'b0101111100100000;
    mem[ 581 ] = 16'b0101111110000001;
    mem[ 582 ] = 16'b0101111111100010;
    mem[ 583 ] = 16'b0110000001000001;
    mem[ 584 ] = 16'b0110000010100001;
    mem[ 585 ] = 16'b0110000011111111;
    mem[ 586 ] = 16'b0110000101011101;
    mem[ 587 ] = 16'b0110000110111001;
    mem[ 588 ] = 16'b0110001000010101;
    mem[ 589 ] = 16'b0110001001110001;
    mem[ 590 ] = 16'b0110001011001011;
    mem[ 591 ] = 16'b0110001100100101;
    mem[ 592 ] = 16'b0110001101111110;
    mem[ 593 ] = 16'b0110001111010110;
    mem[ 594 ] = 16'b0110010000101110;
    mem[ 595 ] = 16'b0110010010000100;
    mem[ 596 ] = 16'b0110010011011010;
    mem[ 597 ] = 16'b0110010100110000;
    mem[ 598 ] = 16'b0110010110000100;
    mem[ 599 ] = 16'b0110010111011000;
    mem[ 600 ] = 16'b0110011000101010;
    mem[ 601 ] = 16'b0110011001111101;
    mem[ 602 ] = 16'b0110011011001110;
    mem[ 603 ] = 16'b0110011100011110;
    mem[ 604 ] = 16'b0110011101101110;
    mem[ 605 ] = 16'b0110011110111101;
    mem[ 606 ] = 16'b0110100000001100;
    mem[ 607 ] = 16'b0110100001011001;
    mem[ 608 ] = 16'b0110100010100110;
    mem[ 609 ] = 16'b0110100011110010;
    mem[ 610 ] = 16'b0110100100111101;
    mem[ 611 ] = 16'b0110100110000111;
    mem[ 612 ] = 16'b0110100111010001;
    mem[ 613 ] = 16'b0110101000011010;
    mem[ 614 ] = 16'b0110101001100010;
    mem[ 615 ] = 16'b0110101010101010;
    mem[ 616 ] = 16'b0110101011110001;
    mem[ 617 ] = 16'b0110101100110111;
    mem[ 618 ] = 16'b0110101101111100;
    mem[ 619 ] = 16'b0110101111000000;
    mem[ 620 ] = 16'b0110110000000100;
    mem[ 621 ] = 16'b0110110001000111;
    mem[ 622 ] = 16'b0110110010001010;
    mem[ 623 ] = 16'b0110110011001011;
    mem[ 624 ] = 16'b0110110100001100;
    mem[ 625 ] = 16'b0110110101001101;
    mem[ 626 ] = 16'b0110110110001100;
    mem[ 627 ] = 16'b0110110111001011;
    mem[ 628 ] = 16'b0110111000001001;
    mem[ 629 ] = 16'b0110111001000110;
    mem[ 630 ] = 16'b0110111010000011;
    mem[ 631 ] = 16'b0110111010111111;
    mem[ 632 ] = 16'b0110111011111011;
    mem[ 633 ] = 16'b0110111100110101;
    mem[ 634 ] = 16'b0110111101101111;
    mem[ 635 ] = 16'b0110111110101001;
    mem[ 636 ] = 16'b0110111111100001;
    mem[ 637 ] = 16'b0111000000011001;
    mem[ 638 ] = 16'b0111000001010001;
    mem[ 639 ] = 16'b0111000010000111;
    mem[ 640 ] = 16'b0111000010111101;
    mem[ 641 ] = 16'b0111000011110011;
    mem[ 642 ] = 16'b0111000100101000;
    mem[ 643 ] = 16'b0111000101011100;
    mem[ 644 ] = 16'b0111000110001111;
    mem[ 645 ] = 16'b0111000111000010;
    mem[ 646 ] = 16'b0111000111110101;
    mem[ 647 ] = 16'b0111001000100110;
    mem[ 648 ] = 16'b0111001001010111;
    mem[ 649 ] = 16'b0111001010001000;
    mem[ 650 ] = 16'b0111001010111000;
    mem[ 651 ] = 16'b0111001011100111;
    mem[ 652 ] = 16'b0111001100010110;
    mem[ 653 ] = 16'b0111001101000100;
    mem[ 654 ] = 16'b0111001101110010;
    mem[ 655 ] = 16'b0111001110011111;
    mem[ 656 ] = 16'b0111001111001011;
    mem[ 657 ] = 16'b0111001111110111;
    mem[ 658 ] = 16'b0111010000100010;
    mem[ 659 ] = 16'b0111010001001101;
    mem[ 660 ] = 16'b0111010001110111;
    mem[ 661 ] = 16'b0111010010100001;
    mem[ 662 ] = 16'b0111010011001010;
    mem[ 663 ] = 16'b0111010011110011;
    mem[ 664 ] = 16'b0111010100011011;
    mem[ 665 ] = 16'b0111010101000011;
    mem[ 666 ] = 16'b0111010101101010;
    mem[ 667 ] = 16'b0111010110010000;
    mem[ 668 ] = 16'b0111010110110110;
    mem[ 669 ] = 16'b0111010111011100;
    mem[ 670 ] = 16'b0111011000000001;
    mem[ 671 ] = 16'b0111011000100110;
    mem[ 672 ] = 16'b0111011001001010;
    mem[ 673 ] = 16'b0111011001101101;
    mem[ 674 ] = 16'b0111011010010001;
    mem[ 675 ] = 16'b0111011010110011;
    mem[ 676 ] = 16'b0111011011010110;
    mem[ 677 ] = 16'b0111011011110111;
    mem[ 678 ] = 16'b0111011100011001;
    mem[ 679 ] = 16'b0111011100111010;
    mem[ 680 ] = 16'b0111011101011010;
    mem[ 681 ] = 16'b0111011101111010;
    mem[ 682 ] = 16'b0111011110011010;
    mem[ 683 ] = 16'b0111011110111001;
    mem[ 684 ] = 16'b0111011111011000;
    mem[ 685 ] = 16'b0111011111110110;
    mem[ 686 ] = 16'b0111100000010100;
    mem[ 687 ] = 16'b0111100000110001;
    mem[ 688 ] = 16'b0111100001001111;
    mem[ 689 ] = 16'b0111100001101011;
    mem[ 690 ] = 16'b0111100010001000;
    mem[ 691 ] = 16'b0111100010100100;
    mem[ 692 ] = 16'b0111100010111111;
    mem[ 693 ] = 16'b0111100011011010;
    mem[ 694 ] = 16'b0111100011110101;
    mem[ 695 ] = 16'b0111100100010000;
    mem[ 696 ] = 16'b0111100100101010;
    mem[ 697 ] = 16'b0111100101000011;
    mem[ 698 ] = 16'b0111100101011101;
    mem[ 699 ] = 16'b0111100101110110;
    mem[ 700 ] = 16'b0111100110001110;
    mem[ 701 ] = 16'b0111100110100111;
    mem[ 702 ] = 16'b0111100110111111;
    mem[ 703 ] = 16'b0111100111010110;
    mem[ 704 ] = 16'b0111100111101101;
    mem[ 705 ] = 16'b0111101000000100;
    mem[ 706 ] = 16'b0111101000011011;
    mem[ 707 ] = 16'b0111101000110001;
    mem[ 708 ] = 16'b0111101001000111;
    mem[ 709 ] = 16'b0111101001011101;
    mem[ 710 ] = 16'b0111101001110010;
    mem[ 711 ] = 16'b0111101010001000;
    mem[ 712 ] = 16'b0111101010011100;
    mem[ 713 ] = 16'b0111101010110001;
    mem[ 714 ] = 16'b0111101011000101;
    mem[ 715 ] = 16'b0111101011011001;
    mem[ 716 ] = 16'b0111101011101101;
    mem[ 717 ] = 16'b0111101100000000;
    mem[ 718 ] = 16'b0111101100010011;
    mem[ 719 ] = 16'b0111101100100110;
    mem[ 720 ] = 16'b0111101100111000;
    mem[ 721 ] = 16'b0111101101001011;
    mem[ 722 ] = 16'b0111101101011101;
    mem[ 723 ] = 16'b0111101101101110;
    mem[ 724 ] = 16'b0111101110000000;
    mem[ 725 ] = 16'b0111101110010001;
    mem[ 726 ] = 16'b0111101110100010;
    mem[ 727 ] = 16'b0111101110110011;
    mem[ 728 ] = 16'b0111101111000011;
    mem[ 729 ] = 16'b0111101111010100;
    mem[ 730 ] = 16'b0111101111100100;
    mem[ 731 ] = 16'b0111101111110011;
    mem[ 732 ] = 16'b0111110000000011;
    mem[ 733 ] = 16'b0111110000010010;
    mem[ 734 ] = 16'b0111110000100001;
    mem[ 735 ] = 16'b0111110000110000;
    mem[ 736 ] = 16'b0111110000111111;
    mem[ 737 ] = 16'b0111110001001101;
    mem[ 738 ] = 16'b0111110001011100;
    mem[ 739 ] = 16'b0111110001101010;
    mem[ 740 ] = 16'b0111110001111000;
    mem[ 741 ] = 16'b0111110010000101;
    mem[ 742 ] = 16'b0111110010010011;
    mem[ 743 ] = 16'b0111110010100000;
    mem[ 744 ] = 16'b0111110010101101;
    mem[ 745 ] = 16'b0111110010111010;
    mem[ 746 ] = 16'b0111110011000110;
    mem[ 747 ] = 16'b0111110011010011;
    mem[ 748 ] = 16'b0111110011011111;
    mem[ 749 ] = 16'b0111110011101011;
    mem[ 750 ] = 16'b0111110011110111;
    mem[ 751 ] = 16'b0111110100000011;
    mem[ 752 ] = 16'b0111110100001111;
    mem[ 753 ] = 16'b0111110100011010;
    mem[ 754 ] = 16'b0111110100100101;
    mem[ 755 ] = 16'b0111110100110000;
    mem[ 756 ] = 16'b0111110100111011;
    mem[ 757 ] = 16'b0111110101000110;
    mem[ 758 ] = 16'b0111110101010001;
    mem[ 759 ] = 16'b0111110101011011;
    mem[ 760 ] = 16'b0111110101100101;
    mem[ 761 ] = 16'b0111110101101111;
    mem[ 762 ] = 16'b0111110101111001;
    mem[ 763 ] = 16'b0111110110000011;
    mem[ 764 ] = 16'b0111110110001101;
    mem[ 765 ] = 16'b0111110110010110;
    mem[ 766 ] = 16'b0111110110100000;
    mem[ 767 ] = 16'b0111110110101001;
    mem[ 768 ] = 16'b0111110110110010;
    mem[ 769 ] = 16'b0111110110111011;
    mem[ 770 ] = 16'b0111110111000100;
    mem[ 771 ] = 16'b0111110111001101;
    mem[ 772 ] = 16'b0111110111010101;
    mem[ 773 ] = 16'b0111110111011110;
    mem[ 774 ] = 16'b0111110111100110;
    mem[ 775 ] = 16'b0111110111101110;
    mem[ 776 ] = 16'b0111110111110110;
    mem[ 777 ] = 16'b0111110111111110;
    mem[ 778 ] = 16'b0111111000000110;
    mem[ 779 ] = 16'b0111111000001110;
    mem[ 780 ] = 16'b0111111000010101;
    mem[ 781 ] = 16'b0111111000011101;
    mem[ 782 ] = 16'b0111111000100100;
    mem[ 783 ] = 16'b0111111000101100;
    mem[ 784 ] = 16'b0111111000110011;
    mem[ 785 ] = 16'b0111111000111010;
    mem[ 786 ] = 16'b0111111001000001;
    mem[ 787 ] = 16'b0111111001000111;
    mem[ 788 ] = 16'b0111111001001110;
    mem[ 789 ] = 16'b0111111001010101;
    mem[ 790 ] = 16'b0111111001011011;
    mem[ 791 ] = 16'b0111111001100010;
    mem[ 792 ] = 16'b0111111001101000;
    mem[ 793 ] = 16'b0111111001101110;
    mem[ 794 ] = 16'b0111111001110101;
    mem[ 795 ] = 16'b0111111001111011;
    mem[ 796 ] = 16'b0111111010000001;
    mem[ 797 ] = 16'b0111111010000110;
    mem[ 798 ] = 16'b0111111010001100;
    mem[ 799 ] = 16'b0111111010010010;
    mem[ 800 ] = 16'b0111111010010111;
    mem[ 801 ] = 16'b0111111010011101;
    mem[ 802 ] = 16'b0111111010100010;
    mem[ 803 ] = 16'b0111111010101000;
    mem[ 804 ] = 16'b0111111010101101;
    mem[ 805 ] = 16'b0111111010110010;
    mem[ 806 ] = 16'b0111111010110111;
    mem[ 807 ] = 16'b0111111010111100;
    mem[ 808 ] = 16'b0111111011000001;
    mem[ 809 ] = 16'b0111111011000110;
    mem[ 810 ] = 16'b0111111011001011;
    mem[ 811 ] = 16'b0111111011010000;
    mem[ 812 ] = 16'b0111111011010100;
    mem[ 813 ] = 16'b0111111011011001;
    mem[ 814 ] = 16'b0111111011011110;
    mem[ 815 ] = 16'b0111111011100010;
    mem[ 816 ] = 16'b0111111011100110;
    mem[ 817 ] = 16'b0111111011101011;
    mem[ 818 ] = 16'b0111111011101111;
    mem[ 819 ] = 16'b0111111011110011;
    mem[ 820 ] = 16'b0111111011110111;
    mem[ 821 ] = 16'b0111111011111011;
    mem[ 822 ] = 16'b0111111011111111;
    mem[ 823 ] = 16'b0111111100000011;
    mem[ 824 ] = 16'b0111111100000111;
    mem[ 825 ] = 16'b0111111100001011;
    mem[ 826 ] = 16'b0111111100001111;
    mem[ 827 ] = 16'b0111111100010010;
    mem[ 828 ] = 16'b0111111100010110;
    mem[ 829 ] = 16'b0111111100011010;
    mem[ 830 ] = 16'b0111111100011101;
    mem[ 831 ] = 16'b0111111100100001;
    mem[ 832 ] = 16'b0111111100100100;
    mem[ 833 ] = 16'b0111111100101000;
    mem[ 834 ] = 16'b0111111100101011;
    mem[ 835 ] = 16'b0111111100101110;
    mem[ 836 ] = 16'b0111111100110001;
    mem[ 837 ] = 16'b0111111100110101;
    mem[ 838 ] = 16'b0111111100111000;
    mem[ 839 ] = 16'b0111111100111011;
    mem[ 840 ] = 16'b0111111100111110;
    mem[ 841 ] = 16'b0111111101000001;
    mem[ 842 ] = 16'b0111111101000100;
    mem[ 843 ] = 16'b0111111101000111;
    mem[ 844 ] = 16'b0111111101001001;
    mem[ 845 ] = 16'b0111111101001100;
    mem[ 846 ] = 16'b0111111101001111;
    mem[ 847 ] = 16'b0111111101010010;
    mem[ 848 ] = 16'b0111111101010100;
    mem[ 849 ] = 16'b0111111101010111;
    mem[ 850 ] = 16'b0111111101011010;
    mem[ 851 ] = 16'b0111111101011100;
    mem[ 852 ] = 16'b0111111101011111;
    mem[ 853 ] = 16'b0111111101100001;
    mem[ 854 ] = 16'b0111111101100100;
    mem[ 855 ] = 16'b0111111101100110;
    mem[ 856 ] = 16'b0111111101101000;
    mem[ 857 ] = 16'b0111111101101011;
    mem[ 858 ] = 16'b0111111101101101;
    mem[ 859 ] = 16'b0111111101101111;
    mem[ 860 ] = 16'b0111111101110010;
    mem[ 861 ] = 16'b0111111101110100;
    mem[ 862 ] = 16'b0111111101110110;
    mem[ 863 ] = 16'b0111111101111000;
    mem[ 864 ] = 16'b0111111101111010;
    mem[ 865 ] = 16'b0111111101111100;
    mem[ 866 ] = 16'b0111111101111110;
    mem[ 867 ] = 16'b0111111110000000;
    mem[ 868 ] = 16'b0111111110000010;
    mem[ 869 ] = 16'b0111111110000100;
    mem[ 870 ] = 16'b0111111110000110;
    mem[ 871 ] = 16'b0111111110001000;
    mem[ 872 ] = 16'b0111111110001010;
    mem[ 873 ] = 16'b0111111110001100;
    mem[ 874 ] = 16'b0111111110001101;
    mem[ 875 ] = 16'b0111111110001111;
    mem[ 876 ] = 16'b0111111110010001;
    mem[ 877 ] = 16'b0111111110010011;
    mem[ 878 ] = 16'b0111111110010100;
    mem[ 879 ] = 16'b0111111110010110;
    mem[ 880 ] = 16'b0111111110011000;
    mem[ 881 ] = 16'b0111111110011001;
    mem[ 882 ] = 16'b0111111110011011;
    mem[ 883 ] = 16'b0111111110011100;
    mem[ 884 ] = 16'b0111111110011110;
    mem[ 885 ] = 16'b0111111110011111;
    mem[ 886 ] = 16'b0111111110100001;
    mem[ 887 ] = 16'b0111111110100010;
    mem[ 888 ] = 16'b0111111110100100;
    mem[ 889 ] = 16'b0111111110100101;
    mem[ 890 ] = 16'b0111111110100111;
    mem[ 891 ] = 16'b0111111110101000;
    mem[ 892 ] = 16'b0111111110101001;
    mem[ 893 ] = 16'b0111111110101011;
    mem[ 894 ] = 16'b0111111110101100;
    mem[ 895 ] = 16'b0111111110101101;
    mem[ 896 ] = 16'b0111111110101110;
    mem[ 897 ] = 16'b0111111110110000;
    mem[ 898 ] = 16'b0111111110110001;
    mem[ 899 ] = 16'b0111111110110010;
    mem[ 900 ] = 16'b0111111110110011;
    mem[ 901 ] = 16'b0111111110110101;
    mem[ 902 ] = 16'b0111111110110110;
    mem[ 903 ] = 16'b0111111110110111;
    mem[ 904 ] = 16'b0111111110111000;
    mem[ 905 ] = 16'b0111111110111001;
    mem[ 906 ] = 16'b0111111110111010;
    mem[ 907 ] = 16'b0111111110111011;
    mem[ 908 ] = 16'b0111111110111100;
    mem[ 909 ] = 16'b0111111110111101;
    mem[ 910 ] = 16'b0111111110111110;
    mem[ 911 ] = 16'b0111111110111111;
    mem[ 912 ] = 16'b0111111111000000;
    mem[ 913 ] = 16'b0111111111000001;
    mem[ 914 ] = 16'b0111111111000010;
    mem[ 915 ] = 16'b0111111111000011;
    mem[ 916 ] = 16'b0111111111000100;
    mem[ 917 ] = 16'b0111111111000101;
    mem[ 918 ] = 16'b0111111111000110;
    mem[ 919 ] = 16'b0111111111000111;
    mem[ 920 ] = 16'b0111111111001000;
    mem[ 921 ] = 16'b0111111111001001;
    mem[ 922 ] = 16'b0111111111001001;
    mem[ 923 ] = 16'b0111111111001010;
    mem[ 924 ] = 16'b0111111111001011;
    mem[ 925 ] = 16'b0111111111001100;
    mem[ 926 ] = 16'b0111111111001101;
    mem[ 927 ] = 16'b0111111111001110;
    mem[ 928 ] = 16'b0111111111001110;
    mem[ 929 ] = 16'b0111111111001111;
    mem[ 930 ] = 16'b0111111111010000;
    mem[ 931 ] = 16'b0111111111010001;
    mem[ 932 ] = 16'b0111111111010001;
    mem[ 933 ] = 16'b0111111111010010;
    mem[ 934 ] = 16'b0111111111010011;
    mem[ 935 ] = 16'b0111111111010011;
    mem[ 936 ] = 16'b0111111111010100;
    mem[ 937 ] = 16'b0111111111010101;
    mem[ 938 ] = 16'b0111111111010101;
    mem[ 939 ] = 16'b0111111111010110;
    mem[ 940 ] = 16'b0111111111010111;
    mem[ 941 ] = 16'b0111111111010111;
    mem[ 942 ] = 16'b0111111111011000;
    mem[ 943 ] = 16'b0111111111011001;
    mem[ 944 ] = 16'b0111111111011001;
    mem[ 945 ] = 16'b0111111111011010;
    mem[ 946 ] = 16'b0111111111011010;
    mem[ 947 ] = 16'b0111111111011011;
    mem[ 948 ] = 16'b0111111111011011;
    mem[ 949 ] = 16'b0111111111011100;
    mem[ 950 ] = 16'b0111111111011101;
    mem[ 951 ] = 16'b0111111111011101;
    mem[ 952 ] = 16'b0111111111011110;
    mem[ 953 ] = 16'b0111111111011110;
    mem[ 954 ] = 16'b0111111111011111;
    mem[ 955 ] = 16'b0111111111011111;
    mem[ 956 ] = 16'b0111111111100000;
    mem[ 957 ] = 16'b0111111111100000;
    mem[ 958 ] = 16'b0111111111100001;
    mem[ 959 ] = 16'b0111111111100001;
    mem[ 960 ] = 16'b0111111111100010;
    mem[ 961 ] = 16'b0111111111100010;
    mem[ 962 ] = 16'b0111111111100011;
    mem[ 963 ] = 16'b0111111111100011;
    mem[ 964 ] = 16'b0111111111100011;
    mem[ 965 ] = 16'b0111111111100100;
    mem[ 966 ] = 16'b0111111111100100;
    mem[ 967 ] = 16'b0111111111100101;
    mem[ 968 ] = 16'b0111111111100101;
    mem[ 969 ] = 16'b0111111111100110;
    mem[ 970 ] = 16'b0111111111100110;
    mem[ 971 ] = 16'b0111111111100110;
    mem[ 972 ] = 16'b0111111111100111;
    mem[ 973 ] = 16'b0111111111100111;
    mem[ 974 ] = 16'b0111111111101000;
    mem[ 975 ] = 16'b0111111111101000;
    mem[ 976 ] = 16'b0111111111101000;
    mem[ 977 ] = 16'b0111111111101001;
    mem[ 978 ] = 16'b0111111111101001;
    mem[ 979 ] = 16'b0111111111101001;
    mem[ 980 ] = 16'b0111111111101010;
    mem[ 981 ] = 16'b0111111111101010;
    mem[ 982 ] = 16'b0111111111101010;
    mem[ 983 ] = 16'b0111111111101011;
    mem[ 984 ] = 16'b0111111111101011;
    mem[ 985 ] = 16'b0111111111101011;
    mem[ 986 ] = 16'b0111111111101100;
    mem[ 987 ] = 16'b0111111111101100;
    mem[ 988 ] = 16'b0111111111101100;
    mem[ 989 ] = 16'b0111111111101101;
    mem[ 990 ] = 16'b0111111111101101;
    mem[ 991 ] = 16'b0111111111101101;
    mem[ 992 ] = 16'b0111111111101101;
    mem[ 993 ] = 16'b0111111111101110;
    mem[ 994 ] = 16'b0111111111101110;
    mem[ 995 ] = 16'b0111111111101110;
    mem[ 996 ] = 16'b0111111111101110;
    mem[ 997 ] = 16'b0111111111101111;
    mem[ 998 ] = 16'b0111111111101111;
    mem[ 999 ] = 16'b0111111111101111;
    mem[ 1000 ] = 16'b0111111111110000;
    mem[ 1001 ] = 16'b0111111111110000;
    mem[ 1002 ] = 16'b0111111111110000;
    mem[ 1003 ] = 16'b0111111111110000;
    mem[ 1004 ] = 16'b0111111111110000;
    mem[ 1005 ] = 16'b0111111111110001;
    mem[ 1006 ] = 16'b0111111111110001;
    mem[ 1007 ] = 16'b0111111111110001;
    mem[ 1008 ] = 16'b0111111111110001;
    mem[ 1009 ] = 16'b0111111111110010;
    mem[ 1010 ] = 16'b0111111111110010;
    mem[ 1011 ] = 16'b0111111111110010;
    mem[ 1012 ] = 16'b0111111111110010;
    mem[ 1013 ] = 16'b0111111111110010;
    mem[ 1014 ] = 16'b0111111111110011;
    mem[ 1015 ] = 16'b0111111111110011;
    mem[ 1016 ] = 16'b0111111111110011;
    mem[ 1017 ] = 16'b0111111111110011;
    mem[ 1018 ] = 16'b0111111111110011;
    mem[ 1019 ] = 16'b0111111111110100;
    mem[ 1020 ] = 16'b0111111111110100;
    mem[ 1021 ] = 16'b0111111111110100;
    mem[ 1022 ] = 16'b0111111111110100;
    mem[ 1023 ] = 16'b0111111111110100;

    end
    
    assign out = mem[y];
    
endmodule
